module ALU(Ain, Bin, ALUop, out, Z);
	input [15:0] Ain, Bin;
	input [1:0] ALUop;
	output [15:0] out;
	output Z;

	reg [15:0] out;
	reg Z;
	
	always @* begin
		
	end

endmodule
